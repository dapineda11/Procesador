library verilog;
use verilog.vl_types.all;
entity SP_vlg_vec_tst is
end SP_vlg_vec_tst;

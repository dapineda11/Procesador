library verilog;
use verilog.vl_types.all;
entity Procesador_vlg_vec_tst is
end Procesador_vlg_vec_tst;

library verilog;
use verilog.vl_types.all;
entity Sistema_vlg_vec_tst is
end Sistema_vlg_vec_tst;
